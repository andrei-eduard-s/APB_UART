`define DATA_SIZE 8
`define PARITY_SIZE 1
`define BAUD_RATE 1
`define STOP_BITS 2